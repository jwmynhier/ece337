/home/ecegrid/a/mg111/ece337/Lab2/source/adder_8bit.sv