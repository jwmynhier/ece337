// $Id: $
// File name:   sensor_b.sv
// Created:     9/1/2016
// Author:      Joseph Mynhier
// Lab Section: 4
// Version:     1.0  Initial Design Entry
// Description: Behavioral Style Sensor Error Detector
