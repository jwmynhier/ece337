// $Id: mg111
// File name:   moore.sv
// Created:     9/15/2016
// Author:      Joseph Mynhier
// Lab Section: 4
// Version:     1.0  Initial Design Entry
// Description: moore model 1101 sequence detector.

module moore
(
	input wire clk,
	input wire n_rst,
	input wire i,
	output reg o
);

endmodule
