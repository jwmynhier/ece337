/home/ecegrid/a/mg111/ece337/Lab2/source/tb_adder_1bit.sv